module ROM (addr,data);
input [31:0] addr;
output [31:0] data;
reg [31:0] data;
localparam ROM_SIZE = 32;
reg [31:0] ROM_DATA[ROM_SIZE-1:0];

always@(*)
	case(addr[7:0])
	  

	  
	  //add test
	  /*
	  0: data<= 32'b00001000000000000000000000000011;
1: data<= 32'b00001000000000000000000000010111;
2: data<= 32'b00001000000000000000000000011011;
3: data<= 32'b00111100000100000100000000000000;
4: data<= 32'b00111100000110001111111111111111;
5: data<= 32'b00100111000110001111111100000000;
6: data<= 32'b00111100000110011111111111111111;
7: data<= 32'b00100111001110011111111100000000;
8: data<= 32'b10101110000000000000000000001000;
9: data<= 32'b10101110000110000000000000000000;
10: data<= 32'b10101110000110010000000000000100;
11: data<= 32'b00100100000010000000000000000011;
12: data<= 32'b10101110000010000000000000001000;
13: data<= 32'b10001110000110000000000000010000;
14: data<= 32'b00000000000110000010000100000010;
15: data<= 32'b00000000000110000111111100000000;
16: data<= 32'b00000000000011110010111100000010;
17: data<= 32'b10101110000110000000000000001100;
18: data<= 32'b00000000100000000101100000100000;
19: data<= 32'b00000000101000000110000000100000;
20: data<= 32'b00000001100010110001000000100000;
21: data<= 32'b00000000000000000000000000100000;
22: data<= 32'b00001000000000000000000000010101;
23: data<= 32'b10101110000000100000000000010100;
24: data<= 32'b00100100000010000000000000000011;
25: data<= 32'b10101110000010000000000000001000;
26: data<= 32'b00000000000000000000000000001000;
27: data<= 32'b00000000000000000000000000100000;
*/
	  
	 0: data<= 32'b00001000000000000000000000000011;
1: data<= 32'b00001000000000000000000000011111;
2: data<= 32'b00001000000000000000000000100011;
3: data<= 32'b00111100000100000100000000000000;
4: data<= 32'b00111100000110001111111111111111;
5: data<= 32'b00100111000110001111111100000000;
6: data<= 32'b00111100000110011111111111111111;
7: data<= 32'b00100111001110011111111100000000;
8: data<= 32'b10101110000000000000000000001000;
9: data<= 32'b10101110000110000000000000000000;
10: data<= 32'b10101110000110010000000000000100;
11: data<= 32'b00100100000010000000000000000011;
12: data<= 32'b10101110000010000000000000001000;
13: data<= 32'b10001110000110000000000000010000;
14: data<= 32'b00000000000110000010000100000010;
15: data<= 32'b00000000000110000111111100000000;
16: data<= 32'b00000000000011110010111100000010;
17: data<= 32'b10101110000110000000000000001100;
18: data<= 32'b00000000100000000101100000100000;
19: data<= 32'b00000000101000000110000000100000;
20: data<= 32'b00000001011011000101000000100010;
21: data<= 32'b00011001010000000000000000000010;
22: data<= 32'b00000001010000000101100000100000;
23: data<= 32'b00001000000000000000000000010100;
24: data<= 32'b00010001011011000000000000000011;
25: data<= 32'b00000001100010110100100000100010;
26: data<= 32'b00000001001000000110000000100000;
27: data<= 32'b00001000000000000000000000010100;
28: data<= 32'b00000001100000000001000000100000;
29: data<= 32'b00000000000000000000000000100000;
30: data<= 32'b00001000000000000000000000011101;
31: data<= 32'b10101110000000100000000000010100;
32: data<= 32'b00100100000010000000000000000011;
33: data<= 32'b10101110000010000000000000001000;
34: data<= 32'b00000000000000000000000000001000;
35: data<= 32'b00000000000000000000000000100000;

	 

		default:	data <= 32'h0800_0000;
	endcase
endmodule